`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:47:31 12/06/2018 
// Design Name: 
// Module Name:    seg_logic 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module seg_logic(
		input wire clk,
		input wire btn,
		output wire [6:0] seg,
		output wire [3:0] an
    );


/*
			case(num_val)
		      0: digit = 7'b1000000;
				1: digit = 7'b1111001;
				2: digit = 7'b0100100;
				3: digit = 7'b0110000;
				4: digit = 7'b0011001;
				5: digit = 7'b0010010;
				6: digit = 7'b0000010;
				7: digit = 7'b1111000;
				8: digit = 7'b0000000;
				9: digit = 7'b0011000;				
		  endcase*/

endmodule
